----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:50:49 01/03/2021 
-- Design Name: 
-- Module Name:    Full_adder_subtractor_128bit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Full_adder_subtractor_128bit is
    Port ( A : in  STD_LOGIC_VECTOR (0 downto 127);
           B : in  STD_LOGIC_VECTOR (0 downto 127);
           Cin : in  STD_LOGIC;
           Output : out  STD_LOGIC_VECTOR (0 downto 128));
end Full_adder_subtractor_128bit;

architecture Behavioral of Full_adder_subtractor_128bit is

begin


end Behavioral;

